module stopwatch (
  input start_stop,
  input reset,
  input clk,
  output [6:0] hex0,
  output [6:0] hex1,
  output [6:0] hex2,
  output [6:0] hex3);


endmodule
